CircuitMaker Text
5.6
Probes: 1
U2_6
Transient Analysis
0 395 79 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 140 10
176 83 1678 999
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 1846 637
9961490 0
0
6 Title:
5 Name:
0
0
0
26
13 Logic Switch~
5 39 224 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D0
-34 0 -20 8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7479 0 0
2
42159.5 3
0
13 Logic Switch~
5 40 175 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D1
-36 0 -22 8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5690 0 0
2
42159.5 2
0
13 Logic Switch~
5 39 127 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D2
-36 1 -22 9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5617 0 0
2
42159.5 1
0
13 Logic Switch~
5 38 76 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D3
-35 1 -21 9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3903 0 0
2
42159.5 0
0
8 Op-Amp5~
219 351 88 0 5 11
0 2 9 4 3 11
0
0 0 848 0
4 OP07
12 4 40 12
2 U2
13 -11 27 -3
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 256 1 0 0 0
1 U
4452 0 0
2
42159.5 13
0
8 Op-Amp5~
219 181 82 0 5 11
0 2 8 6 5 7
0
0 0 848 0
4 OP07
10 7 38 15
2 U1
10 -14 24 -6
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 256 1 0 0 0
1 U
6282 0 0
2
42159.5 12
0
7 Ground~
168 156 102 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7187 0 0
2
42159.5 11
0
7 Ground~
168 319 110 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6866 0 0
2
42159.5 10
0
2 +V
167 351 117 0 1 3
0 3
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7670 0 0
2
42159.5 9
0
2 +V
167 351 65 0 1 3
0 4
0
0 0 53616 0
4 +15V
-14 -13 14 -5
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
951 0 0
2
42159.5 8
0
2 +V
167 250 29 0 1 3
0 10
0
0 0 53616 90
3 +5V
-11 -15 10 -7
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9536 0 0
2
42159.5 7
0
7 Ground~
168 116 281 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5495 0 0
2
42159.5 6
0
2 +V
167 181 108 0 1 3
0 5
0
0 0 53616 180
4 -15V
-12 3 16 11
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8152 0 0
2
42159.5 5
0
2 +V
167 181 59 0 1 3
0 6
0
0 0 53616 0
4 +15V
-13 -13 15 -5
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6223 0 0
2
42159.5 4
0
11 Resistor:A~
219 347 27 0 2 5
0 9 11
0
0 0 880 0
3 10k
-11 -14 10 -6
3 R10
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5441 0 0
2
42159.5 25
0
11 Resistor:A~
219 285 27 0 3 5
0 10 9 1
0
0 0 880 0
3 10k
-11 -14 10 -6
3 R11
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3189 0 0
2
42159.5 24
0
11 Resistor:A~
219 285 82 0 2 5
0 7 9
0
0 0 880 0
3 10k
-11 -14 10 -6
3 R12
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8460 0 0
2
42159.5 23
0
11 Resistor:A~
219 179 29 0 2 5
0 8 7
0
0 0 880 0
6 21.35k
-21 -14 21 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5179 0 0
2
42159.5 22
0
11 Resistor:A~
219 116 250 0 3 5
0 2 16 -1
0
0 0 880 90
3 20k
5 0 26 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3593 0 0
2
42159.5 21
0
11 Resistor:A~
219 116 199 0 2 5
0 16 17
0
0 0 880 90
3 10k
5 0 26 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3928 0 0
2
42159.5 20
0
11 Resistor:A~
219 116 151 0 2 5
0 17 18
0
0 0 880 90
3 10k
5 0 26 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
363 0 0
2
42159.5 19
0
11 Resistor:A~
219 116 101 0 2 5
0 18 8
0
0 0 880 90
3 10k
5 0 26 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8132 0 0
2
42159.5 18
0
11 Resistor:A~
219 70 224 0 2 5
0 12 16
0
0 0 880 0
3 20k
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
65 0 0
2
42159.5 17
0
11 Resistor:A~
219 69 175 0 2 5
0 15 17
0
0 0 880 0
3 20k
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6609 0 0
2
42159.5 16
0
11 Resistor:A~
219 69 127 0 2 5
0 14 18
0
0 0 880 0
3 20k
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8995 0 0
2
42159.5 15
0
11 Resistor:A~
219 69 76 0 2 5
0 13 8
0
0 0 880 0
3 20k
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3918 0 0
2
42159.5 14
0
27
1 1 2 0 0 8336 0 8 5 0 0 3
319 104
319 94
333 94
4 1 3 0 0 4240 0 5 9 0 0 2
351 101
351 102
3 1 4 0 0 4240 0 5 10 0 0 2
351 75
351 74
4 1 5 0 0 4240 0 6 13 0 0 2
181 95
181 93
3 1 6 0 0 4240 0 6 14 0 0 2
181 69
181 68
1 1 2 0 0 16 0 7 6 0 0 3
156 96
156 88
163 88
2 0 7 0 0 8208 0 18 0 0 10 3
197 29
228 29
228 82
1 0 8 0 0 8336 0 18 0 0 9 3
161 29
116 29
116 76
2 0 8 0 0 16 0 6 0 0 24 2
163 76
116 76
5 1 7 0 0 4240 0 6 17 0 0 2
199 82
267 82
1 0 9 0 0 4112 0 15 0 0 12 2
329 27
317 27
2 0 9 0 0 8336 0 16 0 0 13 3
303 27
317 27
317 82
2 2 9 0 0 16 0 17 5 0 0 2
303 82
333 82
1 1 10 0 0 4240 0 11 16 0 0 2
261 27
267 27
2 5 11 0 0 8336 0 15 5 0 0 4
365 27
393 27
393 88
369 88
1 1 12 0 0 4240 0 1 23 0 0 2
51 224
52 224
1 1 13 0 0 4240 0 4 26 0 0 2
50 76
51 76
1 1 14 0 0 16 0 3 25 0 0 2
51 127
51 127
1 1 15 0 0 4240 0 2 24 0 0 2
52 175
51 175
1 1 2 0 0 16 0 12 19 0 0 2
116 275
116 268
2 0 16 0 0 4240 0 23 0 0 27 2
88 224
116 224
2 0 17 0 0 4240 0 24 0 0 26 2
87 175
116 175
2 0 18 0 0 4240 0 25 0 0 25 2
87 127
116 127
2 2 8 0 0 16 0 26 22 0 0 3
87 76
116 76
116 83
2 1 18 0 0 16 0 21 22 0 0 2
116 133
116 119
2 1 17 0 0 16 0 20 21 0 0 2
116 181
116 169
2 1 16 0 0 16 0 19 20 0 0 2
116 232
116 217
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
