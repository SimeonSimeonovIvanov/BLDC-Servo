CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 130 10
176 83 1022 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.309148 0.500000
344 179 457 276
42991634 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 57 295 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21872 0
2 5V
-29 -4 -15 4
0
15 GATE 3,2 ENABLE
-54 -18 51 -10
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8559 0 0
2
42166.8 12
0
13 Logic Switch~
5 57 262 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21872 0
2 5V
-29 -4 -15 4
0
15 GATE 1,4 ENABLE
-54 -18 51 -10
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3674 0 0
2
42166.8 11
0
13 Logic Switch~
5 57 329 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21872 0
2 5V
-29 -4 -15 4
0
11 GATE ENABLE
-40 -18 37 -10
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5697 0 0
2
42166.8 6
0
13 Logic Switch~
5 57 84 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21872 0
2 5V
-29 -4 -15 4
0
9 DIRECTION
-36 -20 27 -12
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3805 0 0
2
42166.8 2
0
13 Logic Switch~
5 249 214 0 1 11
0 14
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5219 0 0
2
42166.8 1
0
13 Logic Switch~
5 57 139 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-29 -4 -15 4
3 OSC
-19 -19 2 -11
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3795 0 0
2
42166.8 0
0
9 2-In AND~
219 414 192 0 3 22
0 7 6 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3637 0 0
2
42166.8 0
0
9 2-In AND~
219 414 102 0 3 22
0 8 6 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3226 0 0
2
42166.8 0
0
9 2-In AND~
219 345 183 0 3 22
0 9 4 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6966 0 0
2
42166.8 0
0
9 2-In AND~
219 341 93 0 3 22
0 10 5 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9796 0 0
2
42166.8 0
0
14 Logic Display~
6 548 64 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 G2H
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5952 0 0
2
42166.8 16
0
14 Logic Display~
6 462 64 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 G1H
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3649 0 0
2
42166.8 15
0
14 Logic Display~
6 548 154 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 G4L
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3716 0 0
2
42166.8 14
0
14 Logic Display~
6 462 154 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 G3L
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4797 0 0
2
42166.8 13
0
5 4013~
219 190 120 0 6 22
0 14 12 15 11 16 10
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 1 0
1 U
4681 0 0
2
42166.8 5
0
5 4013~
219 190 210 0 6 22
0 14 11 15 12 17 9
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 1 0
1 U
9730 0 0
2
42166.8 4
0
10 2-In NAND~
219 111 174 0 3 22
0 12 12 11
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9874 0 0
2
42166.8 3
0
23
1 0 2 0 0 12432 0 13 0 0 4 5
548 172
548 192
511 192
511 102
462 102
1 0 3 0 0 12432 0 11 0 0 3 5
548 82
548 123
499 123
499 192
462 192
1 3 3 0 0 16 0 14 7 0 0 3
462 172
462 192
435 192
1 3 2 0 0 16 0 12 8 0 0 3
462 82
462 102
435 102
1 2 4 0 0 4240 0 1 9 0 0 4
69 295
304 295
304 192
321 192
1 2 5 0 0 4240 0 2 10 0 0 4
69 262
286 262
286 102
317 102
2 0 6 0 0 4112 0 7 0 0 8 2
390 201
379 201
1 2 6 0 0 4240 0 3 8 0 0 4
69 329
379 329
379 111
390 111
1 3 7 0 0 4240 0 7 9 0 0 2
390 183
366 183
1 3 8 0 0 4240 0 8 10 0 0 2
390 93
362 93
6 1 9 0 0 4240 0 16 9 0 0 2
214 174
321 174
6 1 10 0 0 4240 0 15 10 0 0 2
214 84
317 84
3 0 11 0 0 4112 0 17 0 0 23 2
138 174
156 174
2 0 12 0 0 4112 0 17 0 0 22 2
87 183
78 183
1 0 12 0 0 16 0 17 0 0 22 2
87 165
78 165
0 0 13 0 0 16 0 0 0 0 0 2
93 174
93 174
1 0 14 0 0 4112 0 5 0 0 18 2
250 201
250 143
1 1 14 0 0 12432 0 16 15 0 0 6
190 153
190 143
250 143
250 53
190 53
190 63
1 0 15 0 0 4112 0 6 0 0 21 2
69 139
143 139
1 0 12 0 0 16 0 4 0 0 22 2
69 84
78 84
3 3 15 0 0 8336 0 15 16 0 0 4
166 102
143 102
143 192
166 192
2 4 12 0 0 8336 0 15 16 0 0 5
166 84
78 84
78 226
190 226
190 216
4 2 11 0 0 12432 0 15 16 0 0 5
190 126
190 130
156 130
156 174
166 174
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
